library verilog;
use verilog.vl_types.all;
entity Instruction_Decoder_vlg_vec_tst is
end Instruction_Decoder_vlg_vec_tst;
